module time (
    time,
    time2,
    time3,
    time4,
    time5,
    time6,
    time7,
    time8,
    time9，
    dhsajchshanskcjsajf
    dfnisghjc
    avfbgf
    vfgrafgreh
    