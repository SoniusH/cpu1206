`define PC_WIDTH 10
`define DATA_WIDTH 32
`define REG_ADDR_WIDTH 5